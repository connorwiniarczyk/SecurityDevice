module Mock_KeyPadDecoder (
	input clk, reset   // clk and reset
	
);

endmodule